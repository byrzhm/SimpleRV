`ifndef IMM_TYPES
`define IMM_TYPES

`define IMM_TYPE_WIDTH       3

// ***** Immediate types *****
`define IMM_I           3'b000
`define IMM_S           3'b001
`define IMM_B           3'b010
`define IMM_U           3'b011
`define IMM_J           3'b100

`endif