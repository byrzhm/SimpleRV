`define RF_PATH   cpu.RF
`define DMEM_PATH cpu.DMEM
`define IMEM_PATH cpu.IMEM